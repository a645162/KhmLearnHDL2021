module FU(clk,data2,data2,dout1,dout2);
